`timescale 1ns / 1ps

module tmds_tx (
);

encode encode_r ();
encode encode_g ();
encode encode_b ();

endmodule
